`timescale 1ns/1ns
`include "mux16_1.v"
module mux16_1_tb;
reg[0:15]w;
reg[3:0]s;
wire f;
mux16_1 mux(s,w,f);
initial begin
    $dumpfile("mux16_1_tb.vcd");
    $dumpvars(0,mux16_1_tb);
    w=16'b1010000010101011;s=0;#20;
    w=16'b1010000010101011;s=1;#20;
    w=16'b1010000010101011;s=2;#20;
    w=16'b1010000010101011;s=3;#20;
    w=16'b1010000010101011;s=4;#20;
    w=16'b1010000010101011;s=5;#20;
    w=16'b1010000010101011;s=6;#20;
    w=16'b1010000010101011;s=7;#20;
    w=16'b1010000010101011;s=8;#20;
    w=16'b1010000010101011;s=9;#20;
    w=16'b1010000010101011;s=10;#20;
    w=16'b1010000010101011;s=11;#20;
    w=16'b1010000010101011;s=12;#20;
    w=16'b1010000010101011;s=13;#20;
    w=16'b1010000010101011;s=14;#20;
    w=16'b1010000010101011;s=15;#20;
end
endmodule